// This just verifies that sandpiper.vh has been included.
`ifndef SANDPIPER_VH
  !!!ERROR: SandPiper project's sp_<proj>.vh file must include sandpiper.vh.
`endif
