magic
tech sky130A
timestamp 1622920796
<< viali >>
rect 102718 28781 102738 28799
<< metal1 >>
rect 102715 28807 102801 28812
rect 102715 28799 102773 28807
rect 102715 28781 102718 28799
rect 102738 28781 102773 28799
rect 102715 28779 102773 28781
rect 102800 28779 102801 28807
rect 102715 28774 102801 28779
rect 104169 26312 104281 26348
<< via1 >>
rect 102773 28779 102800 28807
<< metal2 >>
rect 102769 28810 102861 28813
rect 102769 28807 102824 28810
rect 102769 28779 102773 28807
rect 102800 28779 102824 28807
rect 102769 28778 102824 28779
rect 102855 28778 102861 28810
rect 102769 28774 102861 28778
rect 101462 28584 101492 28590
<< via2 >>
rect 102824 28778 102855 28810
<< metal3 >>
rect 102875 28816 102931 28819
rect 102819 28814 102931 28816
rect 102819 28810 102884 28814
rect 102819 28778 102824 28810
rect 102855 28778 102884 28810
rect 102919 28778 102931 28814
rect 102819 28774 102931 28778
rect 102875 28773 102931 28774
rect 104169 26312 104281 26348
<< via3 >>
rect 102884 28778 102919 28814
<< mimcapcontact >>
rect 105103 28779 105138 28813
<< metal4 >>
rect 98736 44448 98784 44455
rect 102882 28814 105143 28816
rect 102882 28778 102884 28814
rect 102919 28813 105143 28814
rect 102919 28779 105103 28813
rect 105138 28779 105143 28813
rect 102919 28778 105143 28779
rect 102882 28776 105143 28778
rect 102882 28774 102978 28776
use 10bitdac_layout  10bitdac_layout_0
timestamp 1622920796
transform 1 0 214 0 1 28846
box -214 -28846 102528 27385
use cap_28p  cap_28p_0
timestamp 1616448691
transform 1 0 105249 0 1 26963
box -984 -1226 12410 12449
<< labels >>
rlabel metal3 104180 26326 104180 26326 1 gnd!
flabel locali s 83000 2734 83029 2792 0 FreeSans 40 0 0 0 VREFL
port 27 nsew signal input
flabel locali s 612 55763 641 55811 0 FreeSans 40 0 0 0 VREFH
port 29 nsew signal input
rlabel metal4 103753 28800 103753 28800 1 OUT
port 30 n signal output
flabel locali s 83503 28493 83503 28493 0 FreeSans 40 0 0 0 D[0]
port 35 nsew signal input
flabel locali s 85026 28829 85053 29225 0 FreeSans 40 0 0 0 D[1]
port 37 nsew signal input
flabel locali s 86780 28343 86822 29263 0 FreeSans 40 0 0 0 D[2]
port 39 nsew signal input
flabel locali s 88491 27461 88524 29297 0 FreeSans 40 0 0 0 D[3]
port 41 nsew signal input
flabel locali s 89913 28403 89945 28950 0 FreeSans 40 0 0 0 D[4]
port 44 nsew signal input
flabel locali s 91584 27439 91608 29302 0 FreeSans 40 0 0 0 D[5]
port 46 nsew signal input
flabel locali s 94200 27425 94235 29321 0 FreeSans 40 0 0 0 D[6]
port 48 nsew signal input
flabel locali s 95945 27443 95982 29360 0 FreeSans 40 0 0 0 D[7]
port 50 nsew signal input
flabel locali s 98048 27418 98086 39855 0 FreeSans 40 0 0 0 D[8]
port 52 nsew signal input
flabel locali s 101395 28692 101506 28740 0 FreeSans 40 0 0 0 D[9]
port 54 nsew signal input
rlabel metal2 101476 28587 101476 28587 1 VSSA
port 57 n ground bidirectional
rlabel metal4 98759 44451 98759 44451 1 VDDA
port 58 n power bidirectional
<< properties >>
string LEFclass CORE
<< end >>
